/**************************************************************************************************
	MODULE: Capture_Unit
	PURPOSE: Take in the inputs and write the sample to all ramQueues every cycle, until triggered
	
	INPUTS:
			
	
	OUTPUTS:
	
	INTERNAL:

**************************************************************************************************/