`timescale 100ps / 10ps
`define EOF 32'hFFFF_FFFF 
`define NULL 0

module LA_dig_tb();

	typedef enum logic [1:0] {ReadReg, WriteReg, Dump} Command;
	typedef enum logic [2:0] {ERR, CH1, CH2, CH3, Ch4, Ch5} Channel;
	typedef enum logic [5:0] {TrigCfg_Reg, CH1TrigCfg_Reg, CH2TrigCfg_Reg, CH3TrigCfg_Reg, CH4TrigCfg_Reg, CH5TrigCfg_Reg, decimator_Reg, VIH_Reg, VIL_Reg, matchH_Reg, matchL_Reg, maskH_Reg, maskL_Reg, baud_cntH_Reg, baud_cntL_Reg, trig_posH_Reg, trig_posL_Reg} Register;
	typedef enum logic [2:0] {IDLE, WRITE, READ, RAM, RESP, ERROR} State;
	
	localparam ACK = 8'hA5;
	localparam NCK = 8'hEE;
	
	parameter ENTRIES = 384,	// defaults to 384 for simulation, use 12288 for DE-0 and 384 for sim
		LOG2 = 9;				// Log base 2 of number of entries, use 14 for DE-0 and 9 for sim
	
	//// Interconnects to DUT/support defined as type wire /////
	wire clk400MHz,locked;			// PLL output signals to DUT
	wire clk;						// 100MHz clock generated at this level from clk400MHz
	wire VIH_PWM,VIL_PWM;			// connect to PWM outputs to monitor
	wire CH1L,CH1H,CH2L,CH2H,CH3L;	// channel data inputs from AFE model
	wire CH3H,CH4L,CH4H,CH5L,CH5H;	// channel data inputs from AFE model
	wire RX,TX;						// interface to host
	wire cmd_sent,resp_rdy;			// from master UART, monitored in test bench
	wire [7:0] resp;				// from master UART, reponse received from DUT
	wire tx_prot;					// UART signal for protocol triggering
	wire SS_n,SCLK,MOSI;			// SPI signals for SPI protocol triggering
	wire CH1L_mux,CH1H_mux;         // output of muxing logic for CH1 to enable testing of protocol triggering
	wire CH2L_mux,CH2H_mux;			// output of muxing logic for CH2 to enable testing of protocol triggering
	wire CH3L_mux,CH3H_mux;			// output of muxing logic for CH3 to enable testing of protocol triggering
	
	////// Stimulus is declared as type reg ///////
	reg REF_CLK, RST_n;
	reg [15:0] host_cmd;			// command host is sending to DUT
	reg send_cmd;					// asserted to initiate sending of command
	reg clr_resp_rdy;				// asserted to knock down resp_rdy
	reg [1:0] clk_div;				// counter used to derive 100MHz clk from clk400MHz
	reg strt_tx;					// kick off unit used for protocol triggering
	
	/////////////////////////////////////////////////////////////
	// Channel Dumps can be written to file to aid in testing //
	///////////////////////////////////////////////////////////
	// setup file pointers here if going to do that
	
	///////////////////////////
	// Define command bytes //
	/////////////////////////
	// May or may not want to make some localparams to represent command bytes to LA core
	
	/////////////////////////////////
	localparam UART_triggering = 1'b0;	// set to true if testing UART based triggering
	localparam SPI_triggering = 1'b1;	// set to true if testing SPI based triggering
	
	
	///// Instantiate Analog Front End model (provides stimulus to channels) ///////
	AFE iAFE(.smpl_clk(clk400MHz),.VIH_PWM(VIH_PWM),.VIL_PWM(VIL_PWM),
			.CH1L(CH1L),.CH1H(CH1H),.CH2L(CH2L),.CH2H(CH2H),.CH3L(CH3L),
			.CH3H(CH3H),.CH4L(CH4L),.CH4H(CH4H),.CH5L(CH5L),.CH5H(CH5H));
			
	//// Mux for muxing in protocol triggering for CH1 /////
	assign {CH1H_mux,CH1L_mux} = (UART_triggering) ? {2{tx_prot}} :		// assign to output of UART_tx used to test UART triggering
								(SPI_triggering) ? {2{SS_n}}: 			// assign to output of SPI SS_n if SPI triggering
								{CH1H,CH1L};
	
	//// Mux for muxing in protocol triggering for CH2 /////
	assign {CH2H_mux,CH2L_mux} = (SPI_triggering) ? {2{SCLK}}: 			// assign to output of SPI SCLK if SPI triggering
								{CH2H,CH2L};	
	
	//// Mux for muxing in protocol triggering for CH3 /////
	assign {CH3H_mux,CH3L_mux} = (SPI_triggering) ? {2{MOSI}}: 			// assign to output of SPI MOSI if SPI triggering
								{CH3H,CH3L};					  
		
	////// Instantiate DUT ////////
	LA_dig iDUT(.clk400MHz(clk400MHz),.RST_n(RST_n),.locked(locked),
				.VIH_PWM(VIH_PWM),.VIL_PWM(VIL_PWM),.CH1L(CH1L_mux),.CH1H(CH1H_mux),
				.CH2L(CH2L_mux),.CH2H(CH2H_mux),.CH3L(CH3L_mux),.CH3H(CH3H_mux),.CH4L(CH4L),
				.CH4H(CH4H),.CH5L(CH5L),.CH5H(CH5H),.RX(RX),.TX(TX));
	
	///// Instantiate PLL to provide 400MHz clk from 50MHz ///////
	pll8x iPLL(.ref_clk(REF_CLK),.RST_n(RST_n),.out_clk(clk400MHz),.locked(locked));
	
	///// It is useful to have a 100MHz clock at this level similar //////
	///// to main system clock (clk).  So we will create one        //////
	always @(posedge clk400MHz, negedge locked)
	if (~locked)
		clk_div <= 2'b00;
	else
		clk_div <= clk_div+1;
	assign clk = clk_div[1];
	
	//// Instantiate Master UART (mimics host commands) //////
	UART_comm_mstr iMSTR(.clk(clk), .rst_n(RST_n), .RX(TX), .TX(RX),
						.cmd(host_cmd), .send_cmd(send_cmd),
						.cmd_sent(cmd_sent), .resp_rdy(resp_rdy),
						.resp(resp), .clr_resp_rdy(clr_resp_rdy));
						
	////////////////////////////////////////////////////////////////
	// Instantiate transmitter as source for protocol triggering //
	//////////////////////////////////////////////////////////////
	UART_tx iTX(.clk(clk), .rst_n(RST_n), .tx(tx_prot), .strt_tx(strt_tx),
			.tx_data(8'h96), .tx_done());
						
	////////////////////////////////////////////////////////////////////
	// Instantiate SPI transmitter as source for protocol triggering //
	//////////////////////////////////////////////////////////////////
	SPI_mstr iSPI(.clk(clk),.rst_n(rst_n),.SS_n(SS_n),.SCLK(SCLK),.wrt(strt_tx),.done(done),
				.data_out(16'h6600),.MOSI(MOSI),.pos_edge(1'b0),.width8(1'b1));
	
	initial begin
	//   put your testing code here.
	end
	
	always
	#100 REF_CLK = ~REF_CLK;
	
	///// Perhaps put some basic tasks in a separate file to keep your test bench less cluttered /////
	`include "tb_tasks.sv"
	
	integer file;
	integer r; 
	logic [80*8:1] command; 
	logic [7:0] addr;
	logic [7:0] data; 
	
	initial 
		begin : file_block 
	  
		file = $fopenr("Test1.txt"); 
		if (file == `NULL) 
			disable file_block; 
	  
		while (!$feof(file)) 
			begin 
			r = $fscanf(file, " %s %h %h \n", command, addr, data); 
			case (command) 
			"INIT": 
				$display("READ mem[%h], expect = %h", addr, data); 
			"READ": 
				$display("WRITE mem[%h] = %h", addr, data); 
			default: 
				$display("Unknown command '%0s'", command); 
			endcase 
			end // while not EOF 
	  
		r = $fcloser(file); 
		end // initial 

endmodule	