module Protocol_Trigger_Unit();